

module TestMux2();

endmodule