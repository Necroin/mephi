

module TestEncoder8to3();

endmodule